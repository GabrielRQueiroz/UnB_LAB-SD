-- Universidade de Brasília
-- Laboratório de Sistemas Digitais
-- Autor: Gabriel Roberto de Queiroz
-- Data: 

-- Cabeçalho com breve descrição

-- ************
-- Circuito:
--
-- ************

-- ************ Package ************
-- constantes e bibliotecas
library IEEE;
use IEEE.std_logic_1164.all

-- ************ Entity ************
-- pinos de entrada e saída


-- ************ Architecture ************
-- implementação do projeto


