library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity exp8visto3 is
  port( clock : in STD_LOGIC;
        ligadesliga : in STD_LOGIC;        
        sensorA : in STD_LOGIC;
        sensorB : in STD_LOGIC;
        num7seg : out STD_LOGIC_VECTOR(7 downto 0);
        displays : out STD_LOGIC_VECTOR(3 downto 0) );
end exp8visto3;

architecture exp8visto3_arch of exp8visto3 is
  -- inserir sinais e componentes aqui 
begin

  -- inserir implementacao aqui 

end exp8visto3_arch;





