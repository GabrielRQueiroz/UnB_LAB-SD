library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity exp8visto2 is
  port( clock : in STD_LOGIC;
        reset : in STD_LOGIC;        
        T60 : out STD_LOGIC;
        T20 : out STD_LOGIC;
        T6 : out STD_LOGIC;
        T5 : out STD_LOGIC;
        num7seg : out STD_LOGIC_VECTOR(7 downto 0);
        displays : out STD_LOGIC_VECTOR(3 downto 0) );
end exp8visto2;

architecture exp8visto2_arch of exp8visto2 is
  -- inserir sinais e componentes aqui 
begin

  -- inserir implementacao aqui 

end exp8visto2_arch;



